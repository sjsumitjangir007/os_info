module main

import os

fn main() {
	println('Hello World!')
	println(os.args)
}
